`timescale 1ns/1ps

module synchronous_fifo_tb;
endmodule
